50	2	0	50
150	10000
40	50
40	50
45	68	10
45	70	30
42	66	10
42	68	10
42	65	10
40	66	20
38	68	20
38	70	10
22	85	10
20	85	40
30	50	10
30	52	20
28	52	20
25	50	10
25	52	40
23	55	10
23	52	10
23	55	20
10	40	30
8	40	40
2	40	20
0	40	30
35	30	10
35	32	10
33	32	20
32	30	10
30	30	10
30	32	30
30	35	10
28	30	10
28	35	10
42	15	10
40	5	30
40	15	40
38	5	30
38	15	10
50	30	10
50	40	50
48	30	10
48	40	10
47	35	10
47	40	10
45	35	10
90	35	10
88	30	10
88	35	20
87	30	10
66	55	10
65	55	20
67	85	20
40	69	20
35	66	10
35	69	10
25	85	20
22	75	30
20	80	40
18	75	20
15	75	20
15	80	10
28	55	10
20	50	10
20	55	10
10	35	20
8	45	20
5	35	10
5	45	10
0	45	20
33	35	10
26	32	10
25	30	10
25	35	10
44	5	20
42	10	40
35	5	20
50	35	20
45	30	10
95	30	30
95	35	20
53	30	10
92	30	10
53	35	50
45	65	20
85	25	10
85	35	30
75	55	20
72	55	10
70	58	20
68	60	30
65	60	30
63	58	10
60	55	10
60	60	10
65	85	40
65	82	10
62	80	30
60	80	10
60	85	30
58	75	20
55	80	10
55	85	20
