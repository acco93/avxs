37	2	0	13
100	10000
30	40
30	40
37	52	7
20	26	9
40	30	21
17	63	19
31	62	23
52	33	11
42	41	19
31	32	29
12	42	21
36	16	10
52	41	15
27	23	3
13	13	9
57	58	28
62	42	8
42	57	8
16	57	16
7	38	28
27	68	7
43	67	14
58	48	6
58	27	19
37	69	11
38	46	12
46	10	23
61	33	26
62	63	17
63	69	6
32	22	9
45	35	15
10	17	27
30	15	16
39	10	10
32	39	5
25	32	25
48	28	18
56	37	10
49	49	30
52	64	16
21	47	15
51	21	5
5	25	23
17	33	41
8	52	10
30	48	15
59	15	14
5	6	7
21	10	13
5	64	11
25	55	17
