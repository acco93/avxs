37	2	0	38
100	10000
40	40
40	40
22	22	18
21	45	11
45	35	30
33	34	19
50	50	15
55	45	16
26	59	29
35	51	16
62	24	8
55	34	17
52	26	13
22	53	28
26	29	27
50	40	19
55	50	10
47	66	24
30	60	16
30	50	33
12	17	15
15	14	11
16	19	18
21	48	17
50	30	21
51	42	27
54	38	19
65	27	14
40	60	21
64	4	13
30	20	18
50	70	9
45	42	30
38	33	10
66	8	11
59	5	3
35	60	1
27	24	6
40	37	20
36	26	26
55	20	21
40	66	26
55	65	37
62	35	12
62	57	31
21	36	19
33	44	20
9	56	13
62	48	15
66	14	22
44	13	28
26	13	12
11	28	6
7	43	27
17	64	14
41	46	18
35	16	29
43	26	22
31	76	25
54	10	12
60	15	14
50	15	19
48	21	20
12	38	5
15	56	22
29	39	12
55	57	22
67	41	16
10	70	7
6	25	26
70	64	24
36	6	15
20	30	11
15	5	28
57	72	37
50	4	8
40	20	10
