90	2	0	30
150	10000
10	45
10	45
25	1	25
25	3	7
31	5	13
32	5	6
31	7	14
32	9	5
34	9	11
35	7	5
34	6	15
35	5	15
40	5	13
39	3	12
36	3	18
73	6	13
73	8	18
24	36	12
76	6	17
76	10	4
76	13	7
78	3	12
78	9	13
79	3	8
79	5	16
79	11	15
82	3	6
82	7	5
84	3	11
84	5	10
84	9	3
85	1	7
87	5	2
85	8	4
87	7	4
86	44	14
86	46	12
92	42	10
94	42	11
94	44	7
96	42	5
83	83	11
85	85	12
85	85	14
85	85	10
87	87	8
87	87	16
90	90	19
90	90	5
93	82	17
93	84	7
94	86	14
95	80	17
37	83	17
35	85	14
35	87	16
44	86	7
46	89	13
46	83	9
46	87	11
46	89	35
48	83	5
50	85	28
10	40	12
18	30	11
17	35	10
16	38	8
14	40	11
15	42	21
11	42	4
18	40	15
21	39	16
20	40	4
18	41	16
20	44	7
22	44	10
20	45	11
20	50	11
22	51	7
18	49	9
16	48	11
20	55	12
18	53	7
14	50	8
15	51	6
16	54	5
13	40	7
15	36	8
18	31	11
25	37	13
16	33	7
25	35	4
46	9	19
47	6	17
90	15	9
86	41	18
85	55	17
89	43	20
89	46	14
89	52	16
92	52	9
94	48	13
99	46	4
99	50	21
83	80	13
93	89	16
99	89	13
50	80	13
50	88	7
54	86	3
54	90	10
10	35	7
16	45	9
25	45	17
30	55	12
28	33	12
33	38	13
30	50	7
30	46	11
25	52	10
5	40	20
5	50	13
