12	2	0	38
100	10000
30	40
30	40
37	52	7
17	63	19
52	33	11
31	32	29
52	41	15
27	23	3
13	13	9
32	22	9
10	17	27
32	39	5
25	32	25
56	37	10
49	49	30
52	64	16
20	26	9
40	30	21
21	47	15
31	62	23
51	21	5
42	41	19
5	25	23
12	42	21
36	16	10
17	33	41
57	58	28
62	42	8
42	57	8
16	57	16
8	52	10
7	38	28
27	68	7
30	48	15
43	67	14
58	48	6
58	27	19
37	69	11
38	46	12
46	10	23
61	33	26
62	63	17
63	69	6
45	35	15
59	15	14
5	6	7
21	10	13
5	64	11
30	15	16
39	10	10
25	55	17
48	28	18
