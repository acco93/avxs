75	2	0	25
150	10000
35	35
35	35
41	49	10
35	17	7
55	45	13
15	30	26
25	30	3
20	50	5
10	43	9
55	60	16
30	60	16
50	35	19
30	25	23
15	10	20
10	20	19
5	30	2
45	20	11
45	10	18
65	20	6
35	40	16
41	37	16
40	60	21
31	52	27
35	69	23
53	52	11
65	55	14
20	20	8
40	25	9
42	7	5
11	14	18
6	38	16
8	56	27
13	52	36
47	47	13
49	58	10
37	31	14
63	23	2
53	12	6
32	12	7
36	26	18
21	24	28
17	34	3
12	24	13
24	58	19
27	69	10
56	39	36
37	47	6
37	56	5
47	16	25
44	17	9
46	13	8
49	11	18
49	42	13
53	43	14
61	52	3
57	48	23
56	37	6
55	54	26
15	47	16
14	37	11
11	31	7
16	22	41
4	18	35
28	18	26
26	52	9
26	35	15
31	67	3
15	19	1
22	22	2
18	24	22
26	27	27
25	24	20
22	27	11
25	21	12
19	21	10
20	26	9
18	18	17
55	20	19
20	65	12
30	5	8
20	40	12
15	60	17
45	65	9
55	5	29
65	35	3
45	30	17
64	42	9
63	65	8
2	60	5
5	5	16
60	12	31
24	12	5
23	3	7
2	48	1
6	68	30
27	43	9
57	29	18
15	77	9
62	77	20
49	73	25
67	5	25
57	68	15
