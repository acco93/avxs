37	2	0	113
150	10000
35	35
35	35
35	17	7
25	30	3
10	43	9
30	60	16
45	10	18
64	42	9
35	69	23
63	65	8
20	20	8
5	5	16
11	14	18
6	38	16
57	29	18
21	24	28
17	34	3
27	69	10
56	39	36
37	47	6
53	43	14
57	48	23
56	37	6
22	22	2
19	21	10
20	26	9
20	26	9
36	16	10
17	33	41
62	42	8
7	38	28
27	68	7
58	48	6
37	69	11
38	46	12
46	10	23
5	6	7
25	32	25
56	37	10
41	49	10
55	45	13
55	20	19
15	30	26
20	50	5
55	60	16
20	65	12
50	35	19
30	25	23
15	10	20
30	5	8
10	20	19
5	30	2
20	40	12
15	60	17
45	65	9
45	20	11
55	5	29
65	35	3
65	20	6
45	30	17
35	40	16
41	37	16
40	60	21
31	52	27
53	52	11
65	55	14
2	60	5
60	12	31
40	25	9
42	7	5
24	12	5
23	3	7
2	48	1
8	56	27
13	52	36
6	68	30
47	47	13
49	58	10
27	43	9
37	31	14
63	23	2
53	12	6
32	12	7
36	26	18
12	24	13
24	58	19
15	77	9
62	77	20
49	73	25
67	5	25
37	56	5
57	68	15
47	16	25
44	17	9
46	13	8
49	11	18
49	42	13
61	52	3
55	54	26
15	47	16
14	37	11
11	31	7
16	22	41
4	18	35
28	18	26
26	52	9
26	35	15
31	67	3
15	19	1
18	24	22
26	27	27
25	24	20
22	27	11
25	21	12
18	18	17
37	52	7
49	49	30
52	64	16
40	30	21
21	47	15
17	63	19
31	62	23
52	33	11
51	21	5
42	41	19
31	32	29
5	25	23
12	42	21
52	41	15
27	23	3
13	13	9
57	58	28
42	57	8
16	57	16
8	52	10
30	48	15
43	67	14
58	27	19
61	33	26
62	63	17
63	69	6
32	22	9
45	35	15
59	15	14
10	17	27
21	10	13
5	64	11
30	15	16
39	10	10
32	39	5
25	55	17
48	28	18
