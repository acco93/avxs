149	2	0	50
150	10000
35	35
35	35
41	49	10
35	17	7
55	45	13
55	20	19
15	30	26
25	30	3
20	50	5
10	43	9
55	60	16
30	60	16
20	65	12
50	35	19
10	20	19
15	60	17
45	65	9
45	20	11
45	10	18
65	35	3
35	40	16
64	42	9
31	52	27
35	69	23
53	52	11
63	65	8
20	20	8
5	5	16
60	12	31
40	25	9
24	12	5
11	14	18
6	38	16
8	56	27
47	47	13
37	31	14
57	29	18
63	23	2
53	12	6
36	26	18
21	24	28
17	34	3
24	58	19
27	69	10
56	39	36
37	47	6
47	16	25
44	17	9
46	13	8
49	11	18
49	42	13
53	43	14
57	48	23
56	37	6
55	54	26
14	37	11
11	31	7
16	22	41
26	52	9
26	35	15
15	19	1
22	22	2
18	24	22
26	27	27
25	24	20
22	27	11
25	21	12
19	21	10
20	26	9
18	18	17
37	52	7
49	49	30
52	64	16
20	26	9
40	30	21
21	47	15
17	63	19
31	62	23
52	33	11
51	21	5
31	32	29
12	42	21
36	16	10
52	41	15
27	23	3
17	33	41
13	13	9
57	58	28
62	42	8
16	57	16
7	38	28
27	68	7
30	48	15
43	67	14
58	48	6
58	27	19
37	69	11
38	46	12
46	10	23
61	33	26
62	63	17
45	35	15
59	15	14
5	6	7
10	17	27
32	39	5
25	32	25
25	55	17
48	28	18
56	37	10
22	22	18
36	26	26
21	45	11
45	35	30
55	20	21
33	34	19
50	50	15
55	45	16
26	59	29
40	66	26
55	65	37
35	51	16
62	35	12
62	24	8
9	56	13
44	13	28
26	13	12
11	28	6
7	43	27
17	64	14
41	46	18
55	34	17
35	16	29
43	26	22
26	29	27
50	40	19
55	50	10
54	10	12
60	15	14
47	66	24
30	60	16
30	50	33
12	17	15
15	14	11
16	19	18
21	48	17
50	30	21
51	42	27
50	15	19
48	21	20
12	38	5
30	25	23
15	10	20
30	5	8
5	30	2
20	40	12
55	5	29
65	20	6
45	30	17
41	37	16
40	60	21
65	55	14
2	60	5
42	7	5
23	3	7
2	48	1
13	52	36
6	68	30
49	58	10
27	43	9
32	12	7
12	24	13
15	77	9
62	77	20
49	73	25
67	5	25
37	56	5
57	68	15
61	52	3
15	47	16
4	18	35
28	18	26
31	67	3
42	41	19
5	25	23
42	57	8
8	52	10
63	69	6
32	22	9
21	10	13
5	64	11
30	15	16
39	10	10
62	57	31
21	36	19
33	44	20
62	48	15
66	14	22
52	26	13
31	76	25
22	53	28
