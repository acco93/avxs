50	2	0	50
150	10000
35	35
35	35
41	49	10
55	45	13
15	30	26
25	30	3
30	25	23
10	20	19
45	20	11
45	10	18
65	20	6
35	40	16
40	60	21
35	69	23
53	52	11
20	20	8
40	25	9
42	7	5
37	31	14
63	23	2
53	12	6
36	26	18
21	24	28
17	34	3
12	24	13
27	69	10
56	39	36
37	47	6
47	16	25
44	17	9
46	13	8
49	11	18
49	42	13
53	43	14
57	48	23
56	37	6
55	54	26
14	37	11
11	31	7
16	22	41
28	18	26
31	67	3
15	19	1
22	22	2
18	24	22
26	27	27
25	24	20
22	27	11
25	21	12
19	21	10
20	26	9
18	18	17
35	17	7
55	20	19
20	50	5
10	43	9
55	60	16
30	60	16
20	65	12
50	35	19
15	10	20
30	5	8
5	30	2
20	40	12
15	60	17
45	65	9
55	5	29
65	35	3
45	30	17
41	37	16
64	42	9
31	52	27
65	55	14
63	65	8
2	60	5
5	5	16
60	12	31
24	12	5
23	3	7
11	14	18
6	38	16
2	48	1
8	56	27
13	52	36
6	68	30
47	47	13
49	58	10
27	43	9
57	29	18
32	12	7
24	58	19
15	77	9
62	77	20
49	73	25
67	5	25
37	56	5
57	68	15
61	52	3
15	47	16
4	18	35
26	52	9
26	35	15
